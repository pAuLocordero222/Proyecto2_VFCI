class scoreboard extends uvm?scoreboard;
    

endclass