class driver extends uvm_driver;
    `uvm_component_utils(driver)

    function new (string name = "driver", uvm_component parent = null);
        super.new (name, parent);
    endfunction

    \\Code

endclass